module generated_module(var_0, var_1, var_2, var_3, var_4, x);
    input [12:0] var_0;
    input [12:0] var_1;
    input [13:0] var_2;
    input [13:0] var_3;
    input [7:0] var_4;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8;

    assign constraint_0 = |((~((var_3 << 14'h9))));
    assign constraint_1 = |(((var_2 - 16'h39dd) + 16'he8c3));
    assign constraint_2 = |(((!(var_1)) ^ 1'h1));
    assign constraint_3 = |(((~(var_4)) / 8'h3));
    assign constraint_4 = |(((!(var_0)) >> 1'h0));
    assign constraint_5 = |(((var_2 >> 14'h1) ^ var_1));
    assign constraint_6 = |(((!(var_0)) && var_3));
    assign constraint_7 = |((~(((~(var_4)) * var_4))));
    assign constraint_8 = |(8'h3);

    assign x = constraint_6 & constraint_2 & constraint_4 & constraint_0 & constraint_7 & constraint_5 & constraint_1 & constraint_3 & constraint_8;
endmodule
