module split_7(var_15, x);
    input [4:0] var_15;
    output wire x;

    assign x = 1 || var_15;
endmodule
