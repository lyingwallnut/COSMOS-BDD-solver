module split_11(var_28, x);
        input [10:0] var_28;
    output wire x;

    assign x = 1'b1;
endmodule
