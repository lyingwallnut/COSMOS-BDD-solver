module split_7(var_13, x);
    input [31:0] var_13;
    output wire x;

    wire constraint_13;

    assign constraint_13 = |((!((var_13 + 32'h75f0b4e2))));
    assign x = constraint_13;
endmodule
