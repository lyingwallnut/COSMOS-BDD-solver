module split_14(var_32, x);
    input [9:0] var_32;
    output wire x;

    assign x = 1 || var_32;
endmodule
