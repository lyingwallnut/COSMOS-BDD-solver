module split_5(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [27:0] var_0;
    input [23:0] var_1;
    input [26:0] var_2;
    input [25:0] var_3;
    input [16:0] var_4;
    input [19:0] var_5;
    input [29:0] var_6;
    input [24:0] var_7;
    input [25:0] var_8;
    input [29:0] var_9;
    input [29:0] var_10;
    input [31:0] var_11;
    input [31:0] var_12;
    input [20:0] var_13;
    input [18:0] var_14;
    input [18:0] var_15;
    input [31:0] var_16;
    input [23:0] var_17;
    input [25:0] var_18;
    input [23:0] var_19;
    output wire x;

    wire constraint_1;

    assign constraint_1 = |((var_13 != 32'h12fda3));
    assign x = constraint_1;
endmodule
