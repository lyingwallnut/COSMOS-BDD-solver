module split_10(var_27, x);
        input [8:0] var_27;
    output wire x;

    assign x = 1'b1;
endmodule
