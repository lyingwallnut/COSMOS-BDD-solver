module split_6(var_12, x);
    input [13:0] var_12;
    output wire x;

    wire constraint_6;

    assign constraint_6 = |((var_12 | 14'h2cd9));
    assign x = constraint_6;
endmodule
