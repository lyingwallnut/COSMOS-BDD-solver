module split_4(var_9, x);
    input [7:0] var_9;
    output wire x;

    assign x = 1 || var_9;
endmodule
