module split_2(var_7, var_17, var_24, x);
    input [14:0] var_7;
    input [14:0] var_17;
    input [8:0] var_24;
    output wire x;

    wire constraint_7, constraint_13, constraint_20, constraint_36, constraint_45;

    assign constraint_7 = |(((~(var_7)) + var_17));
    assign constraint_13 = |((~((var_24 - 16'h62))));
    assign constraint_20 = |(((var_17 - 16'h2d49) << 16'hc));
    assign constraint_36 = |(((var_17 || var_24) - 16'h0));
    assign constraint_45 = |((!((var_24 << 9'h0))));
    assign x = constraint_13 & constraint_45 & constraint_36 & constraint_7 & constraint_20;
endmodule
