module split_17(var_38, x);
    input [8:0] var_38;
    output wire x;

    assign x = 1 || var_38;
endmodule
