module split_16(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, var_40, var_41, var_42, var_43, var_44, var_45, var_46, var_47, var_48, var_49, x);
    input [4:0] var_0;
    input [4:0] var_1;
    input [6:0] var_2;
    input [6:0] var_3;
    input [4:0] var_4;
    input [4:0] var_5;
    input [5:0] var_6;
    input [5:0] var_7;
    input [6:0] var_8;
    input [7:0] var_9;
    input [7:0] var_10;
    input [3:0] var_11;
    input [3:0] var_12;
    input [3:0] var_13;
    input [6:0] var_14;
    input [7:0] var_15;
    input [3:0] var_16;
    input [5:0] var_17;
    input [4:0] var_18;
    input [7:0] var_19;
    input [7:0] var_20;
    input [3:0] var_21;
    input [6:0] var_22;
    input [6:0] var_23;
    input [7:0] var_24;
    input [6:0] var_25;
    input [5:0] var_26;
    input [6:0] var_27;
    input [7:0] var_28;
    input [3:0] var_29;
    input [3:0] var_30;
    input [7:0] var_31;
    input [7:0] var_32;
    input [6:0] var_33;
    input [3:0] var_34;
    input [4:0] var_35;
    input [3:0] var_36;
    input [4:0] var_37;
    input [3:0] var_38;
    input [6:0] var_39;
    input [3:0] var_40;
    input [7:0] var_41;
    input [7:0] var_42;
    input [6:0] var_43;
    input [3:0] var_44;
    input [3:0] var_45;
    input [7:0] var_46;
    input [6:0] var_47;
    input [7:0] var_48;
    input [7:0] var_49;
    output wire x;

    assign x = 1'b1;
endmodule
