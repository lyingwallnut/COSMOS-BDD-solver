module split_5(var_15, x);
        input [14:0] var_15;
    output wire x;

    assign x = 1'b1;
endmodule
