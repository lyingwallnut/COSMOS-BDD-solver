module split_21(var_44, x);
    input [14:0] var_44;
    output wire x;

    assign x = 1 || var_44;
endmodule
