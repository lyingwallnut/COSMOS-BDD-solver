module split_12(var_29, x);
        input [12:0] var_29;
    output wire x;

    assign x = 1'b1;
endmodule
