module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, x);
    input [29:0] var_0;
    input [17:0] var_1;
    input [14:0] var_2;
    input [28:0] var_3;
    input [6:0] var_4;
    input [10:0] var_5;
    input [7:0] var_6;
    input [16:0] var_7;
    input [6:0] var_8;
    input [21:0] var_9;
    input [12:0] var_10;
    input [14:0] var_11;
    input [9:0] var_12;
    input [21:0] var_13;
    input [4:0] var_14;
    input [3:0] var_15;
    input [6:0] var_16;
    input [16:0] var_17;
    input [31:0] var_18;
    input [23:0] var_19;
    input [17:0] var_20;
    input [15:0] var_21;
    input [6:0] var_22;
    input [22:0] var_23;
    input [16:0] var_24;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24;

    assign constraint_0 = |(((~(var_17)) && var_7));
    assign constraint_1 = |(((var_19 << 24'h9) != 32'h213a0b));
    assign constraint_2 = |((var_12 - 32'h30a));
    assign constraint_3 = |((var_10 && var_13));
    assign constraint_4 = |((~((var_22 * var_14))));
    assign constraint_5 = |(((var_17 - var_2) >> 17'ha));
    assign constraint_6 = |((!((!((var_24 + var_2))))));
    assign constraint_7 = |(((~(var_24)) + var_12));
    assign constraint_8 = |((var_6 != var_20));
    assign constraint_9 = |(((~(var_11)) + var_1));
    assign constraint_10 = |(((var_24 + var_3) ^ var_7));
    assign constraint_11 = |((var_6 - var_4));
    assign constraint_12 = |((var_22 + 32'h16));
    assign constraint_13 = |((~(((!(var_21)) - 32'h0))));
    assign constraint_14 = |((var_1 || var_19));
    assign constraint_15 = |((var_3 | var_13));
    assign constraint_16 = |((~(((~(var_5)) & var_4))));
    assign constraint_17 = |((!(var_7 != 0) || (var_5 != 0)));
    assign constraint_18 = |(((!(var_16)) != var_3));
    assign constraint_19 = |(((var_15 * 8'hb) ^ var_16));
    assign constraint_20 = |(((!(var_11)) != 32'h1));
    assign constraint_21 = |((var_16 | var_8));
    assign constraint_22 = |((!(((!(var_12)) || var_4))));
    assign constraint_23 = |(((!(var_15)) * var_14));
    assign constraint_24 = |((var_17 ^ 17'h198d3));

    assign x = constraint_21 & constraint_12 & constraint_22 & constraint_11 & constraint_2 & constraint_23 & constraint_16 & constraint_4 & constraint_8 & constraint_3 & constraint_7 & constraint_19 & constraint_0 & constraint_20 & constraint_24 & constraint_9 & constraint_14 & constraint_13 & constraint_6 & constraint_17 & constraint_18 & constraint_5 & constraint_10 & constraint_15 & constraint_1;
endmodule
