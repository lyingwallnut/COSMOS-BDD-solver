module split_1(var_2, x);
    input [10:0] var_2;
    output wire x;

    assign x = 1 || var_2;
endmodule
