module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [27:0] var_0;
    input [23:0] var_1;
    input [26:0] var_2;
    input [25:0] var_3;
    input [16:0] var_4;
    input [19:0] var_5;
    input [29:0] var_6;
    input [24:0] var_7;
    input [25:0] var_8;
    input [29:0] var_9;
    input [29:0] var_10;
    input [31:0] var_11;
    input [31:0] var_12;
    input [20:0] var_13;
    input [18:0] var_14;
    input [18:0] var_15;
    input [31:0] var_16;
    input [23:0] var_17;
    input [25:0] var_18;
    input [23:0] var_19;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19;

    assign constraint_0 = |((var_0 + var_12));
    assign constraint_1 = |((var_13 != 32'h12fda3));
    assign constraint_2 = |((~(((!(var_18)) - var_6))));
    assign constraint_3 = |(((var_19 - var_0) != var_10));
    assign constraint_4 = |(((var_12 || var_9) >> 1'h0));
    assign constraint_5 = |(((var_14 << 19'h4) & var_15));
    assign constraint_6 = |((var_15 && var_2));
    assign constraint_7 = |(((!(var_16)) - var_9));
    assign constraint_8 = |(((var_17 != 32'hd4cb6d) || var_3));
    assign constraint_9 = |(((!(var_8)) || var_17));
    assign constraint_10 = |((var_18 + var_14));
    assign constraint_11 = |((var_0 & 28'hcc7bcd2));
    assign constraint_12 = |((!(((~(var_19)) || var_6))));
    assign constraint_13 = |((var_7 | 25'h3c0e8c));
    assign constraint_14 = |((var_19 & 24'h3fefcb));
    assign constraint_15 = |(((var_8 >> 26'h6) - 32'h3f96300));
    assign constraint_16 = |(((var_0 | var_4) || var_17));
    assign constraint_17 = |(((~(var_4)) + var_8));
    assign constraint_18 = |(((var_14 + var_4) && var_18));
    assign constraint_19 = |((var_8 ^ var_18));

    assign x = constraint_1 & constraint_5 & constraint_18 & constraint_6 & constraint_10 & constraint_17 & constraint_14 & constraint_16 & constraint_9 & constraint_13 & constraint_8 & constraint_11 & constraint_12 & constraint_15 & constraint_19 & constraint_3 & constraint_0 & constraint_2 & constraint_4 & constraint_7;
endmodule
