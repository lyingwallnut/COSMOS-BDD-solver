module split_1(var_5, x);
        input [11:0] var_5;
    output wire x;

    assign x = 1'b1;
endmodule
