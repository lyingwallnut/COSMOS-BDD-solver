module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, var_40, var_41, var_42, var_43, var_44, var_45, var_46, var_47, var_48, var_49, var_50, var_51, var_52, var_53, var_54, var_55, var_56, var_57, var_58, var_59, var_60, var_61, var_62, var_63, var_64, var_65, var_66, var_67, var_68, var_69, var_70, var_71, var_72, var_73, var_74, var_75, var_76, var_77, var_78, var_79, var_80, var_81, var_82, var_83, var_84, var_85, var_86, var_87, var_88, var_89, var_90, var_91, var_92, var_93, var_94, var_95, var_96, var_97, var_98, var_99, var_100, var_101, var_102, var_103, var_104, var_105, var_106, var_107, var_108, var_109, var_110, var_111, var_112, var_113, var_114, var_115, var_116, var_117, var_118, var_119, var_120, var_121, var_122, var_123, var_124, var_125, var_126, var_127, var_128, var_129, var_130, var_131, var_132, var_133, var_134, var_135, var_136, var_137, var_138, var_139, var_140, var_141, var_142, var_143, var_144, var_145, var_146, var_147, var_148, var_149, x);
    input [9:0] var_0;
    input [10:0] var_1;
    input [9:0] var_2;
    input [13:0] var_3;
    input [6:0] var_4;
    input [15:0] var_5;
    input [10:0] var_6;
    input [14:0] var_7;
    input [8:0] var_8;
    input [10:0] var_9;
    input [6:0] var_10;
    input [11:0] var_11;
    input [13:0] var_12;
    input [11:0] var_13;
    input [10:0] var_14;
    input [14:0] var_15;
    input [4:0] var_16;
    input [3:0] var_17;
    input [3:0] var_18;
    input [5:0] var_19;
    input [9:0] var_20;
    input [9:0] var_21;
    input [9:0] var_22;
    input [7:0] var_23;
    input [3:0] var_24;
    input [3:0] var_25;
    input [6:0] var_26;
    input [15:0] var_27;
    input [10:0] var_28;
    input [5:0] var_29;
    input [15:0] var_30;
    input [8:0] var_31;
    input [11:0] var_32;
    input [14:0] var_33;
    input [4:0] var_34;
    input [4:0] var_35;
    input [9:0] var_36;
    input [12:0] var_37;
    input [9:0] var_38;
    input [5:0] var_39;
    input [14:0] var_40;
    input [11:0] var_41;
    input [11:0] var_42;
    input [4:0] var_43;
    input [15:0] var_44;
    input [9:0] var_45;
    input [13:0] var_46;
    input [5:0] var_47;
    input [7:0] var_48;
    input [4:0] var_49;
    input [4:0] var_50;
    input [3:0] var_51;
    input [15:0] var_52;
    input [5:0] var_53;
    input [14:0] var_54;
    input [13:0] var_55;
    input [7:0] var_56;
    input [15:0] var_57;
    input [14:0] var_58;
    input [4:0] var_59;
    input [14:0] var_60;
    input [9:0] var_61;
    input [4:0] var_62;
    input [12:0] var_63;
    input [10:0] var_64;
    input [5:0] var_65;
    input [7:0] var_66;
    input [8:0] var_67;
    input [4:0] var_68;
    input [12:0] var_69;
    input [7:0] var_70;
    input [9:0] var_71;
    input [11:0] var_72;
    input [11:0] var_73;
    input [12:0] var_74;
    input [14:0] var_75;
    input [15:0] var_76;
    input [3:0] var_77;
    input [7:0] var_78;
    input [9:0] var_79;
    input [7:0] var_80;
    input [12:0] var_81;
    input [10:0] var_82;
    input [9:0] var_83;
    input [10:0] var_84;
    input [9:0] var_85;
    input [11:0] var_86;
    input [12:0] var_87;
    input [7:0] var_88;
    input [13:0] var_89;
    input [8:0] var_90;
    input [15:0] var_91;
    input [12:0] var_92;
    input [8:0] var_93;
    input [4:0] var_94;
    input [15:0] var_95;
    input [8:0] var_96;
    input [8:0] var_97;
    input [13:0] var_98;
    input [8:0] var_99;
    input [3:0] var_100;
    input [15:0] var_101;
    input [5:0] var_102;
    input [15:0] var_103;
    input [10:0] var_104;
    input [13:0] var_105;
    input [4:0] var_106;
    input [13:0] var_107;
    input [10:0] var_108;
    input [8:0] var_109;
    input [10:0] var_110;
    input [8:0] var_111;
    input [3:0] var_112;
    input [8:0] var_113;
    input [13:0] var_114;
    input [4:0] var_115;
    input [4:0] var_116;
    input [7:0] var_117;
    input [8:0] var_118;
    input [9:0] var_119;
    input [11:0] var_120;
    input [14:0] var_121;
    input [11:0] var_122;
    input [11:0] var_123;
    input [6:0] var_124;
    input [10:0] var_125;
    input [3:0] var_126;
    input [7:0] var_127;
    input [5:0] var_128;
    input [14:0] var_129;
    input [3:0] var_130;
    input [5:0] var_131;
    input [10:0] var_132;
    input [4:0] var_133;
    input [4:0] var_134;
    input [11:0] var_135;
    input [15:0] var_136;
    input [11:0] var_137;
    input [5:0] var_138;
    input [14:0] var_139;
    input [3:0] var_140;
    input [9:0] var_141;
    input [11:0] var_142;
    input [10:0] var_143;
    input [15:0] var_144;
    input [8:0] var_145;
    input [10:0] var_146;
    input [13:0] var_147;
    input [6:0] var_148;
    input [15:0] var_149;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_27, constraint_28, constraint_29, constraint_30, constraint_31, constraint_32, constraint_33, constraint_34, constraint_35, constraint_36, constraint_37, constraint_38, constraint_39, constraint_40, constraint_41, constraint_42, constraint_43, constraint_44, constraint_45, constraint_46, constraint_47, constraint_48, constraint_49, constraint_50, constraint_51, constraint_52, constraint_53, constraint_54, constraint_55, constraint_56, constraint_57, constraint_58, constraint_59, constraint_60, constraint_61, constraint_62, constraint_63, constraint_64, constraint_65, constraint_66, constraint_67, constraint_68, constraint_69, constraint_70, constraint_71, constraint_72, constraint_73, constraint_74, constraint_75, constraint_76, constraint_77, constraint_78, constraint_79, constraint_80, constraint_81, constraint_82, constraint_83, constraint_84, constraint_85, constraint_86, constraint_87, constraint_88, constraint_89, constraint_90, constraint_91, constraint_92, constraint_93, constraint_94, constraint_95, constraint_96, constraint_97, constraint_98, constraint_99, constraint_100, constraint_101, constraint_102, constraint_103, constraint_104;

    assign constraint_0 = |((var_31 & var_26));
    assign constraint_1 = |(((-var_62) ^ var_77));
    assign constraint_2 = |(((~(var_24)) & var_17));
    assign constraint_3 = |((var_141 >> 10'h0));
    assign constraint_4 = |(((~(var_115)) || var_73));
    assign constraint_5 = |(((var_120 | var_13) && var_110));
    assign constraint_6 = |((var_126 * 8'h9));
    assign constraint_7 = |(((!(var_28)) + 16'h1));
    assign constraint_8 = |(((~(var_102)) - 16'h3d));
    assign constraint_9 = |(((~(var_46)) && var_85));
    assign constraint_10 = |(((-var_125) && var_67));
    assign constraint_11 = |((!(var_10 != 0) || (var_34 != 0)));
    assign constraint_12 = |(((~(var_22)) || var_91));
    assign constraint_13 = |((var_39 - var_143));
    assign constraint_14 = |(((-var_108) << 11'h2));
    assign constraint_15 = |(((-var_85) | var_71));
    assign constraint_16 = |(((var_128 ^ var_62) != 16'h30));
    assign constraint_17 = |(((-var_140) / 4'h5));
    assign constraint_18 = |((var_59 != 16'h17));
    assign constraint_19 = |(((~(var_135)) >> 12'h8));
    assign constraint_20 = |((var_126 && var_66));
    assign constraint_21 = |(((var_138 ^ 6'h18) >> 6'h0));
    assign constraint_22 = |(((!(var_70)) - var_116));
    assign constraint_23 = |((var_20 << 10'h5));
    assign constraint_24 = |((var_51 / 4'h8));
    assign constraint_25 = |(((var_27 || var_82) - var_58));
    assign constraint_26 = |(((-var_145) ^ var_67));
    assign constraint_27 = |(((var_2 + var_35) || var_55));
    assign constraint_28 = |((var_71 & 10'h2a9));
    assign constraint_29 = |((var_117 + var_42));
    assign constraint_30 = |(((-var_67) - 16'h1d1));
    assign constraint_31 = |(((!(var_12)) >> 1'h0));
    assign constraint_32 = |((var_111 || var_20));
    assign constraint_33 = |((var_69 >> 13'h9));
    assign constraint_34 = |((var_108 - 16'h40b));
    assign constraint_35 = |(((!(var_129)) || var_72));
    assign constraint_36 = |(((var_113 << 9'h7) | var_127));
    assign constraint_37 = |((var_148 != var_61));
    assign constraint_38 = |(((var_73 & var_49) << 12'h0));
    assign constraint_39 = |((var_31 << 9'h2));
    assign constraint_40 = |(((!(var_144)) << 1'h0));
    assign constraint_41 = |(((~(var_81)) && var_81));
    assign constraint_42 = |((!((~(var_51)) != 0) || (4'h2 != 0)));
    assign constraint_43 = |(((~(var_0)) && var_31));
    assign constraint_44 = |((var_8 | 9'h4));
    assign constraint_45 = |(((!(var_87)) || var_88));
    assign constraint_46 = |((var_43 || var_93));
    assign constraint_47 = |((var_137 && var_26));
    assign constraint_48 = |((!((-var_34) != 0) || (5'h7 != 0)));
    assign constraint_49 = |(((var_132 - var_46) & var_142));
    assign constraint_50 = |(((var_44 - 16'he03e) ^ var_86));
    assign constraint_51 = |(((~(var_131)) * 8'h5));
    assign constraint_52 = |(((!(var_144)) != var_12));
    assign constraint_53 = |((var_131 && var_78));
    assign constraint_54 = |(((!(var_124)) << 1'h0));
    assign constraint_55 = |((var_2 + 16'h12b));
    assign constraint_56 = |(((var_48 >> 8'h1) >> 8'h2));
    assign constraint_57 = |(((var_5 & var_75) >> 16'hb));
    assign constraint_58 = |(((var_92 ^ var_50) & var_51));
    assign constraint_59 = |((var_78 / 8'hf));
    assign constraint_60 = |(((var_125 - 16'h6b8) || var_78));
    assign constraint_61 = |((var_133 + var_112));
    assign constraint_62 = |(((-var_46) || var_123));
    assign constraint_63 = |(((var_33 ^ var_19) ^ var_135));
    assign constraint_64 = |(((var_115 | 5'h1e) || var_116));
    assign constraint_65 = |(((-var_123) - var_2));
    assign constraint_66 = |((var_52 || var_38));
    assign constraint_67 = |(((!(var_108)) != 16'h1));
    assign constraint_68 = |(((var_77 / 4'hb) + 16'hc));
    assign constraint_69 = |(((var_33 - 16'h6e36) + 16'hdf10));
    assign constraint_70 = |(((~(var_117)) - var_33));
    assign constraint_71 = |((var_19 ^ 6'h3d));
    assign constraint_72 = |((var_53 || var_79));
    assign constraint_73 = |((var_148 & var_77));
    assign constraint_74 = |((var_54 - 16'h1bde));
    assign constraint_75 = |((var_15 & var_115));
    assign constraint_76 = |(((var_140 && var_11) != 16'h0));
    assign constraint_77 = |(((var_112 / 4'h2) ^ var_18));
    assign constraint_78 = |(((-var_104) >> 11'h2));
    assign constraint_79 = |((var_10 * 8'hb));
    assign constraint_80 = |(((var_37 << 13'h4) ^ var_111));
    assign constraint_81 = |(((-var_46) ^ var_80));
    assign constraint_82 = |(((var_31 ^ 9'h10d) || var_17));
    assign constraint_83 = |((var_138 != var_84));
    assign constraint_84 = |(((var_66 >> 8'h2) ^ 8'ha7));
    assign constraint_85 = |(((var_144 << 16'h6) | 16'h8622));
    assign constraint_86 = |((var_99 << 9'h4));
    assign constraint_87 = |((var_38 & 10'h9e));
    assign constraint_88 = |(((~(var_0)) ^ var_83));
    assign constraint_89 = |((var_44 & var_33));
    assign constraint_90 = |((var_146 ^ var_96));
    assign constraint_91 = |(((!(var_112)) * var_51));
    assign constraint_92 = |(((var_94 * var_117) << 8'h1));
    assign constraint_93 = |((!((~(var_81)) != 0) || (var_41 != 0)));
    assign constraint_94 = |(((var_51 + var_62) | 5'h8));
    assign constraint_95 = |((var_66 || var_39));
    assign constraint_96 = |(((var_18 != 16'h0) + var_71));
    assign constraint_97 = |((!((-var_122) != 0) || (var_65 != 0)));
    assign constraint_98 = |((var_5 + var_95));
    assign constraint_99 = |(((var_11 + 16'hba9) >> 16'h4));
    assign constraint_100 = |(4'h2);
    assign constraint_101 = |(4'h5);
    assign constraint_102 = |(4'h8);
    assign constraint_103 = |(4'hb);
    assign constraint_104 = |(8'hf);

    assign x = constraint_61 & constraint_18 & constraint_2 & constraint_20 & constraint_73 & constraint_95 & constraint_53 & constraint_64 & constraint_46 & constraint_42 & constraint_94 & constraint_8 & constraint_11 & constraint_72 & constraint_22 & constraint_48 & constraint_54 & constraint_0 & constraint_71 & constraint_6 & constraint_13 & constraint_83 & constraint_47 & constraint_4 & constraint_37 & constraint_32 & constraint_1 & constraint_39 & constraint_86 & constraint_91 & constraint_44 & constraint_76 & constraint_96 & constraint_16 & constraint_82 & constraint_43 & constraint_55 & constraint_23 & constraint_56 & constraint_87 & constraint_21 & constraint_28 & constraint_75 & constraint_29 & constraint_3 & constraint_60 & constraint_38 & constraint_45 & constraint_36 & constraint_27 & constraint_30 & constraint_10 & constraint_51 & constraint_79 & constraint_34 & constraint_58 & constraint_90 & constraint_7 & constraint_97 & constraint_9 & constraint_15 & constraint_84 & constraint_66 & constraint_67 & constraint_92 & constraint_70 & constraint_5 & constraint_78 & constraint_65 & constraint_12 & constraint_14 & constraint_88 & constraint_19 & constraint_26 & constraint_41 & constraint_33 & constraint_35 & constraint_99 & constraint_62 & constraint_49 & constraint_93 & constraint_74 & constraint_80 & constraint_81 & constraint_25 & constraint_31 & constraint_89 & constraint_52 & constraint_98 & constraint_63 & constraint_40 & constraint_69 & constraint_57 & constraint_50 & constraint_85 & constraint_24 & constraint_68 & constraint_17 & constraint_59 & constraint_77 & constraint_100 & constraint_101 & constraint_102 & constraint_103 & constraint_104;
endmodule
