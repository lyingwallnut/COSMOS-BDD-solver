module split_13(var_30, x);
        input [6:0] var_30;
    output wire x;

    assign x = 1'b1;
endmodule
