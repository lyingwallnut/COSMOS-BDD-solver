module split_8(var_18, x);
    input [8:0] var_18;
    output wire x;

    assign x = 1 || var_18;
endmodule
