module split_9(var_19, x);
    input [28:0] var_19;
    output wire x;

    assign x = 1 || var_19;
endmodule
