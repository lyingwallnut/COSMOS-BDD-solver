module split_5(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [26:0] var_0;
    input [40:0] var_1;
    input [28:0] var_2;
    input [51:0] var_3;
    input [45:0] var_4;
    input [24:0] var_5;
    input [16:0] var_6;
    input [28:0] var_7;
    input [5:0] var_8;
    input [37:0] var_9;
    input [46:0] var_10;
    input [40:0] var_11;
    input [26:0] var_12;
    input [51:0] var_13;
    input [26:0] var_14;
    input [39:0] var_15;
    input [28:0] var_16;
    input [52:0] var_17;
    input [7:0] var_18;
    input [19:0] var_19;
    output wire x;

    assign x = 1'b1;
endmodule
