module split_11(var_23, x);
    input [11:0] var_23;
    output wire x;

    assign x = 1 || var_23;
endmodule
