module split_8(var_17, x);
    input [28:0] var_17;
    output wire x;

    assign x = 1 || var_17;
endmodule
