module split_0(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, var_40, var_41, var_42, var_43, var_44, var_45, var_46, var_47, var_48, var_49, x);
    input [10:0] var_0;
    input [3:0] var_1;
    input [10:0] var_2;
    input [5:0] var_3;
    input [11:0] var_4;
    input [11:0] var_5;
    input [4:0] var_6;
    input [14:0] var_7;
    input [12:0] var_8;
    input [7:0] var_9;
    input [3:0] var_10;
    input [5:0] var_11;
    input [4:0] var_12;
    input [14:0] var_13;
    input [15:0] var_14;
    input [4:0] var_15;
    input [11:0] var_16;
    input [14:0] var_17;
    input [8:0] var_18;
    input [9:0] var_19;
    input [7:0] var_20;
    input [15:0] var_21;
    input [6:0] var_22;
    input [11:0] var_23;
    input [8:0] var_24;
    input [9:0] var_25;
    input [14:0] var_26;
    input [12:0] var_27;
    input [10:0] var_28;
    input [3:0] var_29;
    input [9:0] var_30;
    input [14:0] var_31;
    input [9:0] var_32;
    input [14:0] var_33;
    input [3:0] var_34;
    input [13:0] var_35;
    input [5:0] var_36;
    input [12:0] var_37;
    input [8:0] var_38;
    input [5:0] var_39;
    input [13:0] var_40;
    input [8:0] var_41;
    input [15:0] var_42;
    input [13:0] var_43;
    input [14:0] var_44;
    input [15:0] var_45;
    input [3:0] var_46;
    input [5:0] var_47;
    input [4:0] var_48;
    input [15:0] var_49;
    output wire x;

    wire constraint_0, constraint_1, constraint_3, constraint_4, constraint_5, constraint_6, constraint_9, constraint_10, constraint_11, constraint_12, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_21, constraint_24, constraint_25, constraint_26, constraint_28, constraint_29, constraint_30, constraint_31, constraint_32, constraint_34, constraint_35, constraint_37, constraint_38, constraint_39, constraint_40, constraint_42, constraint_43, constraint_44, constraint_47, constraint_48, constraint_49, constraint_50, constraint_51, constraint_52;

    assign constraint_0 = |(((var_36 / 6'hd) + var_0));
    assign constraint_1 = |(((~(var_5)) | var_10));
    assign constraint_3 = |((~(((~(var_27)) && var_22))));
    assign constraint_4 = |((~(((~(var_26)) >> 15'h5))));
    assign constraint_5 = |((!((var_12 * var_3) != 0) || (6'h26 != 0)));
    assign constraint_6 = |((var_29 & 4'h8));
    assign constraint_9 = |(((~(var_10)) << 4'h1));
    assign constraint_10 = |((var_10 ^ 4'hc));
    assign constraint_11 = |((var_26 ^ var_22));
    assign constraint_12 = |(((var_36 * 8'h8) & 8'h22));
    assign constraint_14 = |((var_21 != var_10));
    assign constraint_15 = |((var_6 != 16'h1a));
    assign constraint_16 = |((~((~((var_5 | 12'hac3))))));
    assign constraint_17 = |((var_42 || var_1));
    assign constraint_18 = |(((~(var_46)) && var_6));
    assign constraint_19 = |((var_31 ^ var_4));
    assign constraint_21 = |((var_45 || var_29));
    assign constraint_24 = |(((var_36 / 6'h4) || var_0));
    assign constraint_25 = |((var_5 + var_42));
    assign constraint_26 = |(((var_39 ^ var_6) * var_11));
    assign constraint_28 = |((~(((~(var_21)) ^ var_45))));
    assign constraint_29 = |(((var_12 * var_34) & var_29));
    assign constraint_30 = |((var_47 * 8'h2));
    assign constraint_31 = |(((~(var_46)) - 16'he));
    assign constraint_32 = |(((var_26 - 16'h7ca9) - 16'h286b));
    assign constraint_34 = |((!(((!(var_16)) || var_1))));
    assign constraint_35 = |((var_0 + var_10));
    assign constraint_37 = |(((var_34 | var_1) && var_25));
    assign constraint_38 = |((!((~(var_16)) != 0) || (var_46 != 0)));
    assign constraint_39 = |((!((var_22 && var_4))));
    assign constraint_40 = |(((var_47 | var_6) / 6'hb));
    assign constraint_42 = |((var_6 && var_27));
    assign constraint_43 = |(((var_39 | 6'h2c) - 16'h39));
    assign constraint_44 = |((var_21 & var_22));
    assign constraint_47 = |(((var_5 >> 12'h3) + 16'h60a));
    assign constraint_48 = |((var_45 || var_29));
    assign constraint_49 = |(((~(var_47)) << 6'h3));
    assign constraint_50 = |(6'h4);
    assign constraint_51 = |(6'hb);
    assign constraint_52 = |(6'hd);
    assign x = constraint_6 & constraint_18 & constraint_15 & constraint_31 & constraint_9 & constraint_10 & constraint_49 & constraint_37 & constraint_35 & constraint_42 & constraint_43 & constraint_1 & constraint_34 & constraint_21 & constraint_48 & constraint_17 & constraint_39 & constraint_14 & constraint_38 & constraint_30 & constraint_29 & constraint_3 & constraint_44 & constraint_12 & constraint_5 & constraint_11 & constraint_26 & constraint_47 & constraint_16 & constraint_25 & constraint_19 & constraint_32 & constraint_4 & constraint_28 & constraint_40 & constraint_24 & constraint_0 & constraint_50 & constraint_51 & constraint_52;
endmodule
