module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [47:0] var_0;
    input [53:0] var_1;
    input [20:0] var_2;
    input [5:0] var_3;
    input [5:0] var_4;
    input [16:0] var_5;
    input [63:0] var_6;
    input [5:0] var_7;
    input [38:0] var_8;
    input [54:0] var_9;
    input [57:0] var_10;
    input [53:0] var_11;
    input [31:0] var_12;
    input [61:0] var_13;
    input [46:0] var_14;
    input [36:0] var_15;
    input [42:0] var_16;
    input [37:0] var_17;
    input [27:0] var_18;
    input [63:0] var_19;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21;

    assign constraint_0 = |(((var_3 / 6'he) * var_7));
    assign constraint_1 = |((var_17 != 64'h34d5a910c));
    assign constraint_2 = |((var_3 - 32'h3b));
    assign constraint_3 = |((var_7 + var_18));
    assign constraint_4 = |((var_6 != var_11));
    assign constraint_5 = |((!((var_15 || var_1) != 0) || (1'h0 != 0)));
    assign constraint_6 = |((!(((!(var_2)) - var_4))));
    assign constraint_7 = |((var_18 + var_4));
    assign constraint_8 = |((~(((~(var_3)) * var_4))));
    assign constraint_9 = |((var_6 | var_9));
    assign constraint_10 = |((var_18 != 64'h5b18a6a));
    assign constraint_11 = |((!(var_11 != 0) || (54'h19e5256ac506f0 != 0)));
    assign constraint_12 = |(((!(var_1 != 0) || (54'h2f9a14264d3a30 != 0)) ^ 1'h0));
    assign constraint_13 = |((!((var_3 + 32'h1b) != 0) || (var_2 != 0)));
    assign constraint_14 = |((~(((!(var_5)) - var_3))));
    assign constraint_15 = |((~((var_7 != var_2))));
    assign constraint_16 = |(((var_11 << 54'h11) & var_0));
    assign constraint_17 = |(((~(var_2)) + var_12));
    assign constraint_18 = |((var_12 | 32'h26058782));
    assign constraint_19 = |((var_3 / 6'hc));
    assign constraint_20 = |(6'hc);
    assign constraint_21 = |(6'he);

    assign x = constraint_2 & constraint_8 & constraint_14 & constraint_15 & constraint_6 & constraint_13 & constraint_3 & constraint_7 & constraint_17 & constraint_10 & constraint_18 & constraint_1 & constraint_5 & constraint_16 & constraint_11 & constraint_12 & constraint_4 & constraint_9 & constraint_19 & constraint_0 & constraint_20 & constraint_21;
endmodule
