module split_8(var_25, x);
        input [12:0] var_25;
    output wire x;

    assign x = 1'b1;
endmodule
