module split_77(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, var_40, var_41, var_42, var_43, var_44, var_45, var_46, var_47, var_48, var_49, var_50, var_51, var_52, var_53, var_54, var_55, var_56, var_57, var_58, var_59, var_60, var_61, var_62, var_63, var_64, var_65, var_66, var_67, var_68, var_69, var_70, var_71, var_72, var_73, var_74, var_75, var_76, var_77, var_78, var_79, var_80, var_81, var_82, var_83, var_84, var_85, var_86, var_87, var_88, var_89, var_90, var_91, var_92, var_93, var_94, var_95, var_96, var_97, var_98, var_99, var_100, var_101, var_102, var_103, var_104, var_105, var_106, var_107, var_108, var_109, var_110, var_111, var_112, var_113, var_114, var_115, var_116, var_117, var_118, var_119, var_120, var_121, var_122, var_123, var_124, var_125, var_126, var_127, var_128, var_129, var_130, var_131, var_132, var_133, var_134, var_135, var_136, var_137, var_138, var_139, var_140, var_141, var_142, var_143, var_144, var_145, var_146, var_147, var_148, var_149, x);
    input [9:0] var_0;
    input [10:0] var_1;
    input [9:0] var_2;
    input [13:0] var_3;
    input [6:0] var_4;
    input [15:0] var_5;
    input [10:0] var_6;
    input [14:0] var_7;
    input [8:0] var_8;
    input [10:0] var_9;
    input [6:0] var_10;
    input [11:0] var_11;
    input [13:0] var_12;
    input [11:0] var_13;
    input [10:0] var_14;
    input [14:0] var_15;
    input [4:0] var_16;
    input [3:0] var_17;
    input [3:0] var_18;
    input [5:0] var_19;
    input [9:0] var_20;
    input [9:0] var_21;
    input [9:0] var_22;
    input [7:0] var_23;
    input [3:0] var_24;
    input [3:0] var_25;
    input [6:0] var_26;
    input [15:0] var_27;
    input [10:0] var_28;
    input [5:0] var_29;
    input [15:0] var_30;
    input [8:0] var_31;
    input [11:0] var_32;
    input [14:0] var_33;
    input [4:0] var_34;
    input [4:0] var_35;
    input [9:0] var_36;
    input [12:0] var_37;
    input [9:0] var_38;
    input [5:0] var_39;
    input [14:0] var_40;
    input [11:0] var_41;
    input [11:0] var_42;
    input [4:0] var_43;
    input [15:0] var_44;
    input [9:0] var_45;
    input [13:0] var_46;
    input [5:0] var_47;
    input [7:0] var_48;
    input [4:0] var_49;
    input [4:0] var_50;
    input [3:0] var_51;
    input [15:0] var_52;
    input [5:0] var_53;
    input [14:0] var_54;
    input [13:0] var_55;
    input [7:0] var_56;
    input [15:0] var_57;
    input [14:0] var_58;
    input [4:0] var_59;
    input [14:0] var_60;
    input [9:0] var_61;
    input [4:0] var_62;
    input [12:0] var_63;
    input [10:0] var_64;
    input [5:0] var_65;
    input [7:0] var_66;
    input [8:0] var_67;
    input [4:0] var_68;
    input [12:0] var_69;
    input [7:0] var_70;
    input [9:0] var_71;
    input [11:0] var_72;
    input [11:0] var_73;
    input [12:0] var_74;
    input [14:0] var_75;
    input [15:0] var_76;
    input [3:0] var_77;
    input [7:0] var_78;
    input [9:0] var_79;
    input [7:0] var_80;
    input [12:0] var_81;
    input [10:0] var_82;
    input [9:0] var_83;
    input [10:0] var_84;
    input [9:0] var_85;
    input [11:0] var_86;
    input [12:0] var_87;
    input [7:0] var_88;
    input [13:0] var_89;
    input [8:0] var_90;
    input [15:0] var_91;
    input [12:0] var_92;
    input [8:0] var_93;
    input [4:0] var_94;
    input [15:0] var_95;
    input [8:0] var_96;
    input [8:0] var_97;
    input [13:0] var_98;
    input [8:0] var_99;
    input [3:0] var_100;
    input [15:0] var_101;
    input [5:0] var_102;
    input [15:0] var_103;
    input [10:0] var_104;
    input [13:0] var_105;
    input [4:0] var_106;
    input [13:0] var_107;
    input [10:0] var_108;
    input [8:0] var_109;
    input [10:0] var_110;
    input [8:0] var_111;
    input [3:0] var_112;
    input [8:0] var_113;
    input [13:0] var_114;
    input [4:0] var_115;
    input [4:0] var_116;
    input [7:0] var_117;
    input [8:0] var_118;
    input [9:0] var_119;
    input [11:0] var_120;
    input [14:0] var_121;
    input [11:0] var_122;
    input [11:0] var_123;
    input [6:0] var_124;
    input [10:0] var_125;
    input [3:0] var_126;
    input [7:0] var_127;
    input [5:0] var_128;
    input [14:0] var_129;
    input [3:0] var_130;
    input [5:0] var_131;
    input [10:0] var_132;
    input [4:0] var_133;
    input [4:0] var_134;
    input [11:0] var_135;
    input [15:0] var_136;
    input [11:0] var_137;
    input [5:0] var_138;
    input [14:0] var_139;
    input [3:0] var_140;
    input [9:0] var_141;
    input [11:0] var_142;
    input [10:0] var_143;
    input [15:0] var_144;
    input [8:0] var_145;
    input [10:0] var_146;
    input [13:0] var_147;
    input [6:0] var_148;
    input [15:0] var_149;
    output wire x;

    assign x = 1'b1;
endmodule
