module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [26:0] var_0;
    input [40:0] var_1;
    input [28:0] var_2;
    input [51:0] var_3;
    input [45:0] var_4;
    input [24:0] var_5;
    input [16:0] var_6;
    input [28:0] var_7;
    input [5:0] var_8;
    input [37:0] var_9;
    input [46:0] var_10;
    input [40:0] var_11;
    input [26:0] var_12;
    input [51:0] var_13;
    input [26:0] var_14;
    input [39:0] var_15;
    input [28:0] var_16;
    input [52:0] var_17;
    input [7:0] var_18;
    input [19:0] var_19;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19;

    assign constraint_0 = |(((var_2 + 32'h214c87d) ^ var_6));
    assign constraint_1 = |(((var_0 << 27'h12) >> 27'h3));
    assign constraint_2 = |(((!(var_18)) * var_8));
    assign constraint_3 = |((!((!(var_0)) != 0) || (1'h0 != 0)));
    assign constraint_4 = |((var_5 - var_18));
    assign constraint_5 = |((var_4 != var_6));
    assign constraint_6 = |((!(var_17 != 0) || (var_7 != 0)));
    assign constraint_7 = |(((var_15 >> 40'h9) | 40'ha71ca2ef72));
    assign constraint_8 = |(((var_18 | 8'h4) * 8'ha));
    assign constraint_9 = |((var_14 >> 27'h4));
    assign constraint_10 = |((var_16 + var_12));
    assign constraint_11 = |(((var_2 | var_5) != 64'h1b4e37e1));
    assign constraint_12 = |((var_0 + var_12));
    assign constraint_13 = |(((~(var_7)) + var_14));
    assign constraint_14 = |((var_6 != 64'h608d));
    assign constraint_15 = |(((!(var_6)) + var_0));
    assign constraint_16 = |((var_4 != var_7));
    assign constraint_17 = |((var_1 != 64'h18e69585ec5));
    assign constraint_18 = |(((var_19 && var_7) != 64'h1));
    assign constraint_19 = |(((var_12 != 64'h44a702e) != var_18));

    assign x = constraint_2 & constraint_8 & constraint_4 & constraint_14 & constraint_19 & constraint_15 & constraint_18 & constraint_12 & constraint_9 & constraint_0 & constraint_10 & constraint_11 & constraint_13 & constraint_3 & constraint_1 & constraint_5 & constraint_16 & constraint_17 & constraint_7 & constraint_6;
endmodule
