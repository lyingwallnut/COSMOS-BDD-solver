module split_0(var_0, var_1, var_3, var_4, var_6, var_7, var_8, var_14, var_15, var_16, var_18, var_20, var_21, var_22, var_24, var_25, var_26, var_28, var_29, x);
    input [28:0] var_0;
    input [26:0] var_1;
    input [23:0] var_3;
    input [3:0] var_4;
    input [9:0] var_6;
    input [16:0] var_7;
    input [11:0] var_8;
    input [7:0] var_14;
    input [17:0] var_15;
    input [7:0] var_16;
    input [17:0] var_18;
    input [8:0] var_20;
    input [17:0] var_21;
    input [10:0] var_22;
    input [6:0] var_24;
    input [29:0] var_25;
    input [26:0] var_26;
    input [26:0] var_28;
    input [6:0] var_29;
    output wire x;

    wire constraint_0, constraint_3, constraint_4, constraint_5, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_15, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_28, constraint_29, constraint_30, constraint_31;

    assign constraint_0 = |((var_14 * var_29));
    assign constraint_3 = |((!(var_24 != 0) || (var_29 != 0)));
    assign constraint_4 = |((var_0 || var_3));
    assign constraint_5 = |(((var_7 & var_4) != var_18));
    assign constraint_7 = |((var_28 - var_14));
    assign constraint_8 = |((!(var_21 != 0) || (var_4 != 0)));
    assign constraint_9 = |(((~(var_25)) | var_1));
    assign constraint_10 = |(((var_16 / 8'h4) && var_6));
    assign constraint_11 = |(((var_16 * var_14) != var_21));
    assign constraint_12 = |((!((var_0 + var_26))));
    assign constraint_15 = |(((var_22 + 32'h41e) - 32'h276a248e));
    assign constraint_17 = |((var_26 != var_15));
    assign constraint_18 = |((~((var_21 && var_25))));
    assign constraint_19 = |((!((~((var_24 * 8'h5))))));
    assign constraint_20 = |(((~(var_21)) << 18'h1));
    assign constraint_21 = |((var_26 << 27'h6));
    assign constraint_22 = |((var_20 | var_24));
    assign constraint_23 = |(((!(var_8)) || var_29));
    assign constraint_24 = |((var_21 << 18'h0));
    assign constraint_25 = |((var_25 || var_6));
    assign constraint_26 = |((!((var_4 + var_26))));
    assign constraint_28 = |(((var_1 | var_22) | var_16));
    assign constraint_29 = |((var_14 != 32'hb8));
    assign constraint_30 = |(4'h7);
    assign constraint_31 = |(8'h4);
    assign x = constraint_29 & constraint_3 & constraint_22 & constraint_23 & constraint_0 & constraint_8 & constraint_15 & constraint_19 & constraint_5 & constraint_26 & constraint_28 & constraint_11 & constraint_7 & constraint_24 & constraint_25 & constraint_20 & constraint_17 & constraint_18 & constraint_4 & constraint_21 & constraint_12 & constraint_9 & constraint_10 & constraint_30 & constraint_31;
endmodule
