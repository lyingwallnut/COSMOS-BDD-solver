module split_4(var_10, x);
    input [31:0] var_10;
    output wire x;

    assign x = 1 || var_10;
endmodule
