module split_2(var_5, x);
    input [26:0] var_5;
    output wire x;

    assign x = 1 || var_5;
endmodule
