module split_11(var_27, x);
    input [6:0] var_27;
    output wire x;

    assign x = 1 || var_27;
endmodule
