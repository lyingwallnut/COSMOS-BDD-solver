module split_10(var_20, x);
    input [7:0] var_20;
    output wire x;

    assign x = 1 || var_20;
endmodule
