module split_2(var_8, x);
        input [9:0] var_8;
    output wire x;

    assign x = 1'b1;
endmodule
