module split_5(var_13, x);
    input [14:0] var_13;
    output wire x;

    assign x = 1 || var_13;
endmodule
