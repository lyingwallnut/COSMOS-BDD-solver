module split_18(var_40, x);
    input [13:0] var_40;
    output wire x;

    assign x = 1 || var_40;
endmodule
