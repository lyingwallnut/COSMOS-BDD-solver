module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [47:0] var_0;
    input [53:0] var_1;
    input [20:0] var_2;
    input [5:0] var_3;
    input [5:0] var_4;
    input [16:0] var_5;
    input [63:0] var_6;
    input [5:0] var_7;
    input [38:0] var_8;
    input [54:0] var_9;
    input [57:0] var_10;
    input [53:0] var_11;
    input [31:0] var_12;
    input [61:0] var_13;
    input [46:0] var_14;
    input [36:0] var_15;
    input [42:0] var_16;
    input [37:0] var_17;
    input [27:0] var_18;
    input [63:0] var_19;
    output wire x;

    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20;

    assign constraint_0 = |((var_4 ^ 6'h31));
    assign constraint_1 = |(((var_19 && var_16) & 1'h1));
    assign constraint_2 = |(((!(var_5)) << 1'h0));
    assign constraint_3 = |((~(((!(var_3)) << 1'h0))));
    assign constraint_4 = |((var_0 >> 48'h1b));
    assign constraint_5 = |(((~(var_10)) || var_8));
    assign constraint_6 = |((var_12 + 32'h2aa55980));
    assign constraint_7 = |(((~(var_14)) ^ 47'h7efe2535ca95));
    assign constraint_8 = |(((!(var_4)) / 1'h1));
    assign constraint_9 = |((~((var_7 * 8'hb))));
    assign constraint_10 = |(((~(var_11)) ^ var_0));
    assign constraint_11 = |((var_7 | 6'h14));
    assign constraint_12 = |(((~(var_5)) - 32'h15266));
    assign constraint_13 = |((var_3 + var_12));
    assign constraint_14 = |((var_11 || var_8));
    assign constraint_15 = |(((~(var_19)) || var_15));
    assign constraint_16 = |(((var_9 << 55'h12) ^ var_15));
    assign constraint_17 = |(((var_7 + 8'h4) * 8'h7));
    assign constraint_18 = |((~((var_4 * var_3))));
    assign constraint_19 = |(((var_18 - 32'hd5a2661) && var_13));
    assign constraint_20 = |(1'h1);

    assign x = constraint_11 & constraint_0 & constraint_3 & constraint_9 & constraint_18 & constraint_17 & constraint_2 & constraint_12 & constraint_13 & constraint_6 & constraint_14 & constraint_19 & constraint_4 & constraint_5 & constraint_7 & constraint_16 & constraint_15 & constraint_10 & constraint_1 & constraint_8 & constraint_20;
endmodule
